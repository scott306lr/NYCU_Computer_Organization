/***************************************************
Student Name: ������ �I�a��
Student ID: 0816137 0716241
***************************************************/

`timescale 1ns/1ps

module Ander(
    	input  src1_i,
	input   src2_i,
	output  sum_o
	);
    
/* Write your code HERE */
assign sum_o=src1_i&src2_i;

endmodule